library verilog;
use verilog.vl_types.all;
entity calculadora_main_vlg_vec_tst is
end calculadora_main_vlg_vec_tst;
