library verilog;
use verilog.vl_types.all;
entity calculadora_2_vlg_vec_tst is
end calculadora_2_vlg_vec_tst;
